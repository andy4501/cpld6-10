LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY UP_COUNTER is
PORT( CLK: IN STD_LOGIC;
Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END UP_COUNTER;
ARCHITECTURE a OF UP_COUNTER IS
SIGNAL QN : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL SN : STD_LOGIC;
BEGIN
PROCESS (CLK)
BEGIN
IF CLK'event AND CLK='1' THEN
	IF SN='0' THEN
		IF QN="00010001" THEN
			SN<='1';
		ELSE
			QN<=QN+1;
		END IF;
	ELSE
		QN<="00000000";
		SN<='0';
	END IF;
END IF;
END PROCESS;
Q<=QN;
END a;